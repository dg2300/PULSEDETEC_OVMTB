package pd_pkg;

	import ovm_pkg::*;

	`include "ovm_macros.svh"
	`include "pd_transaction.sv"
    `include "pd_sequencer.sv"
	`include "pd_driver.sv"
	`include "pd_agent.sv"
	`include "pd_env.sv"
	`include "pd_sequence.sv"
	`include "pd_test.sv"

endpackage