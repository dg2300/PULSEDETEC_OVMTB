interface dut_interface;
	logic clock;
	logic reset;
	logic sig_in,sig_out;
	time delay;
endinterface